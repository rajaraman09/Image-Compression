// barrel48
//`include "mux48to1.v"

module barrel48(o,i,s);
input [47:0] i;
input [7:0] s;
output [47:0] o;
wire a;
assign a=1'b0;

mux48to1 mu1(o[0],i[0],i[1],i[2],i[3],i[4],i[5],i[6],i[7],i[8],i[9],i[10],i[11],i[12],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu2(o[1],i[1],i[2],i[3],i[4],i[5],i[6],i[7],i[8],i[9],i[10],i[11],i[12],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu3(o[2],i[2],i[3],i[4],i[5],i[6],i[7],i[8],i[9],i[10],i[11],i[12],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu4(o[3],i[3],i[4],i[5],i[6],i[7],i[8],i[9],i[10],i[11],i[12],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu5(o[4],i[4],i[5],i[6],i[7],i[8],i[9],i[10],i[11],i[12],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu6(o[5],i[5],i[6],i[7],i[8],i[9],i[10],i[11],i[12],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu7(o[6],i[6],i[7],i[8],i[9],i[10],i[11],i[12],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu8(o[7],i[7],i[8],i[9],i[10],i[11],i[12],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu9(o[8],i[8],i[9],i[10],i[11],i[12],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu10(o[9],i[9],i[10],i[11],i[12],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu11(o[10],i[10],i[11],i[12],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu12(o[11],i[11],i[12],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu13(o[12],i[12],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu14(o[13],i[13],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu15(o[14],i[14],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu16(o[15],i[15],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu17(o[16],i[16],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu18(o[17],i[17],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu19(o[18],i[18],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu20(o[19],i[19],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu21(o[20],i[20],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu22(o[21],i[21],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu23(o[22],i[22],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu24(o[23],i[23],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu25(o[24],i[24],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu26(o[25],i[25],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu27(o[26],i[26],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu28(o[27],i[27],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu29(o[28],i[28],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu30(o[29],i[29],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu31(o[30],i[30],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu32(o[31],i[31],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu33(o[32],i[32],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu34(o[33],i[33],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu35(o[34],i[34],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu36(o[35],i[35],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu37(o[36],i[36],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu38(o[37],i[37],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu39(o[38],i[38],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu40(o[39],i[39],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu41(o[40],i[40],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu42(o[41],i[41],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu43(o[42],i[42],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu44(o[43],i[43],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu45(o[44],i[44],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu46(o[45],i[45],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu47(o[46],i[46],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);
mux48to1 mu48(o[47],i[47],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[7],s[6],s[5],s[4],s[3],s[2],s[1],s[0]);

endmodule








































