// barrel 24 bit shifter - left
//`include "mux24to1.v"

module barrel24(o,i,s);
input [23:0] i;
input [4:0] s;
output [23:0] o;
wire a;
assign a=1'b0;

mux24to1 mu1(o[0],i[0],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu2(o[1],i[1],i[0],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu3(o[2],i[2],i[1],i[0],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu4(o[3],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu5(o[4],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu6(o[5],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu7(o[6],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu8(o[7],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu9(o[8],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu10(o[9],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu11(o[10],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu12(o[11],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu13(o[12],i[12],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu14(o[13],i[13],i[12],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu15(o[14],i[14],i[13],i[12],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu16(o[15],i[15],i[14],i[13],i[12],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu17(o[16],i[16],i[15],i[14],i[13],i[12],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu18(o[17],i[17],i[16],i[15],i[14],i[13],i[12],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu19(o[18],i[18],i[17],i[16],i[15],i[14],i[13],i[12],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu20(o[19],i[19],i[18],i[17],i[16],i[15],i[14],i[13],i[12],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu21(o[20],i[20],i[19],i[18],i[17],i[16],i[15],i[14],i[13],i[12],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu22(o[21],i[21],i[20],i[19],i[18],i[17],i[16],i[15],i[14],i[13],i[12],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu23(o[22],i[22],i[21],i[20],i[19],i[18],i[17],i[16],i[15],i[14],i[13],i[12],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],a,s[4],s[3],s[2],s[1],s[0]);
mux24to1 mu24(o[23],i[23],i[22],i[21],i[20],i[19],i[18],i[17],i[16],i[15],i[14],i[13],i[12],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0],s[4],s[3],s[2],s[1],s[0]);

endmodule
