module increment_unsigned_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_1_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_1_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_1_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_10_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_10_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_10_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_11_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_11_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_11_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_12_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_12_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_12_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_13_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_13_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_13_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_14_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_14_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_14_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_15_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_15_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_15_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_16_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_16_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_16_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_17_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_17_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_17_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_18_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_18_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_18_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_19_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_19_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_19_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_2_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_2_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_2_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_20_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_20_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_20_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_21_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_21_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_21_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_22_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_22_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_22_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_23_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_23_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_23_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_24_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_24_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_24_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_25_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_25_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_25_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_26_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_26_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_26_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_27_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_27_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_27_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_28_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_28_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_28_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_29_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_29_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_29_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_3_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_3_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_3_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_30_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_30_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_30_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_31_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_31_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_31_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_32_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_32_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_32_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_33_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_33_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_33_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_34_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_34_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_34_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_35_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_35_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_35_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_36_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_36_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_36_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_37_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_37_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_37_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_38_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_38_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_38_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_39_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_39_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_39_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_4_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_4_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_4_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_40_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_40_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_40_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_41_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_41_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_41_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_42_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_42_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_42_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_43_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_43_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_43_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_44_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_44_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_44_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_45_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_45_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_45_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_46_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_46_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_46_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_47_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_47_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_47_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_5_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_5_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_5_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_6_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_6_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_6_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_7_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_7_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_7_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_8_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_8_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_8_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_9_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_50, A[0], CI);
  xor g24 (Z[1], A[1], n_50);
  and g25 (n_51, A[1], n_50);
  xor g26 (Z[2], A[2], n_51);
  and g27 (n_52, A[2], n_51);
  xor g28 (Z[3], A[3], n_52);
  and g29 (n_53, A[3], n_52);
  xor g30 (Z[4], A[4], n_53);
  and g31 (n_54, A[4], n_53);
  xor g32 (Z[5], A[5], n_54);
  and g33 (n_55, A[5], n_54);
  xor g34 (Z[6], A[6], n_55);
  and g35 (n_56, A[6], n_55);
  xor g36 (Z[7], A[7], n_56);
  and g37 (n_57, A[7], n_56);
  xor g38 (Z[8], A[8], n_57);
  and g39 (n_58, A[8], n_57);
  xor g40 (Z[9], A[9], n_58);
  and g41 (n_59, A[9], n_58);
  xor g42 (Z[10], A[10], n_59);
  and g43 (n_60, A[10], n_59);
  xor g44 (Z[11], A[11], n_60);
  and g45 (n_61, A[11], n_60);
  xor g46 (Z[12], A[12], n_61);
  and g47 (n_62, A[12], n_61);
  xor g48 (Z[13], A[13], n_62);
  and g49 (n_63, A[13], n_62);
  xor g50 (Z[14], A[14], n_63);
  and g51 (n_64, A[14], n_63);
  xor g52 (Z[15], A[15], n_64);
  and g53 (n_65, A[15], n_64);
  xor g54 (Z[16], A[16], n_65);
  and g55 (n_66, A[16], n_65);
  xor g56 (Z[17], A[17], n_66);
  and g57 (n_67, A[17], n_66);
  xor g58 (Z[18], A[18], n_67);
  and g59 (n_68, A[18], n_67);
  xor g60 (Z[19], A[19], n_68);
  and g61 (n_69, A[19], n_68);
  xor g62 (Z[20], A[20], n_69);
  and g63 (n_70, A[20], n_69);
  xor g64 (Z[21], A[21], n_70);
  and g65 (n_71, A[21], n_70);
  xor g66 (Z[22], A[22], n_71);
  and g67 (n_72, A[22], n_71);
  xor g68 (Z[23], A[23], n_72);
endmodule

module increment_unsigned_9_GENERIC(A, CI, Z);
  input [23:0] A;
  input CI;
  output [23:0] Z;
  wire [23:0] A;
  wire CI;
  wire [23:0] Z;
  increment_unsigned_9_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

